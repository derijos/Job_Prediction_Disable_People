���      �sklearn.preprocessing._label��LabelEncoder���)��}�(�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK'��h	�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�13 years of experience in acute healthcare setting��ASN��	B.Com/BBA��B.E./B.Tech��B.Ed in Education��BSN��)Baccalaureate degree in Nursing or higher��Bachelor in Sonography��Bachelor's degree in psychology��Bachelors Degree��Bachelors Degree in Finance��Bachelors degree in Accounting��Chemical Engineering��Communication��Computer Science��D Pharma��Dental��Diploma in Domestic Plumbing��!Diploma in Electrical Engineering��Doctoral��English Language��GED��HR Analytics��HSE��High School Diploma��Hindi/English Language��M.D./M.S. in Medicine��MBBS��MD��MSN��Masters��Masters in Library Science��Other��PG��!PG degree in financial management��PMP certification��UG��UG/PG��UG/PG in Management�et�b�_sklearn_version��0.23.2�ub.