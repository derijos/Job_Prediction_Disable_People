��b      �numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK'��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�High School Diploma��Bachelors Degree��Chemical Engineering��B.E./B.Tech��Dental��MD��BSN��MBBS��English Language��Computer Science��ASN��PMP certification��Bachelors Degree in Finance��UG/PG��UG/PG in Management��UG��Doctoral��B.Ed in Education��Bachelor's degree in psychology��HSE��!PG degree in financial management��13 years of experience in acute healthcare setting��MSN��Communication��PG��GED��!Diploma in Electrical Engineering��Masters in Library Science��Bachelors degree in Accounting��	B.Com/BBA��D Pharma��)Baccalaureate degree in Nursing or higher��Bachelor in Sonography��Other��Diploma in Domestic Plumbing��Masters��M.D./M.S. in Medicine��Hindi/English Language��HR Analytics�et�b.