�cnumpy.core.multiarray
_reconstruct
q cnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   O8qK K�q	Rq
(KX   |qNNNJ����J����K?tqb�]q(X   2000 - 6999qX   7000 - 14999qX   15000 - 34999qX   35000 - 50000qetqb.