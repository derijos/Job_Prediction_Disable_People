��%      �sklearn.preprocessing._label��LabelEncoder���)��}�(�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h	�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�15000 - 34999��2000 - 6999��35000 - 50000��7000 - 14999�et�b�_sklearn_version��0.23.2�ub.